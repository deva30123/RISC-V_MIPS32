module decode(
  input[31:0] NPC,
  input[31:0] IR,
  input[31:0] rb_in
  output [31:0] A,
  output [31:0] B;
);
  reg [31:0] reg [31:0];
  
endmodule
