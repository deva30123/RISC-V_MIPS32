module inst_mem (
  input write,
  input addr_w,
  input addr_r,
  output read,
)
  
