module decode(
  input[31:0] NPC,
  input[31:0] IR,
  output [31:0] A,
  output [31:0] B;
);
  reg [31:0] reg [31:0];
  
endmodule
