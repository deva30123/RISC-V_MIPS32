module ifetch(
  input ALU,
  input sel,
  output NPC,
  output IR
);
  reg [9:0] PC;
  PC = 
endmodule
